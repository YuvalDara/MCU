-- Ifetch module (provides the PC and instruction memory for the MIPS computer)
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
LIBRARY altera_mf;
USE altera_mf.altera_mf_components.all;


ENTITY Ifetch IS
	generic(
		WORD_GRANULARITY 	: boolean := False;
		DATA_BUS_WIDTH 		: integer := 32;
		PC_WIDTH 				: integer := 10;
		NEXT_PC_WIDTH 		: integer := 8; -- NEXT_PC_WIDTH = PC_WIDTH-2
		ITCM_ADDR_WIDTH 		: integer := 8;
		WORDS_NUM 			: integer := 256;
		INST_CNT_WIDTH 		: integer := 16
	);
	PORT(	
		clk_i, rst_i 		: IN STD_LOGIC;
		add_result_i 		: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        Branch_ctrl_i 	: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		Jump_ctrl_i 		: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		alu_res_i			: IN STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
        zero_i 			: IN STD_LOGIC;
		jump_PC_to_ISR_i : IN STD_LOGIC;
		ISR_addr_i 		: IN STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
		pc_o 			: OUT STD_LOGIC_VECTOR(PC_WIDTH-1 DOWNTO 0);
		pc_plus4_o 		: OUT STD_LOGIC_VECTOR(PC_WIDTH-1 DOWNTO 0);
		instruction_o 	: OUT STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
		inst_cnt_o 		: OUT STD_LOGIC_VECTOR(INST_CNT_WIDTH-1 DOWNTO 0);
		next_pc_no_INT_o	: OUT STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0)
	);
END Ifetch;


ARCHITECTURE behavior OF Ifetch IS
	SIGNAL pc_q				  		: STD_LOGIC_VECTOR(PC_WIDTH-1 DOWNTO 0);
	SIGNAL pc_plus4_r 				: STD_LOGIC_VECTOR(PC_WIDTH-1 DOWNTO 0);
	SIGNAL itcm_addr_w 				: STD_LOGIC_VECTOR(ITCM_ADDR_WIDTH-1 DOWNTO 0);
	SIGNAL next_pc_mux1_w  		: STD_LOGIC_VECTOR(NEXT_PC_WIDTH-1 DOWNTO 0);
	SIGNAL next_pc_mux2_w  		: STD_LOGIC_VECTOR(NEXT_PC_WIDTH-1 DOWNTO 0);
	SIGNAL next_pc_with_interrupts_w 	: STD_LOGIC_VECTOR(NEXT_PC_WIDTH-1 DOWNTO 0);
	SIGNAL rst_flag_q				: STD_LOGIC;
	SIGNAL inst_cnt_q 				: STD_LOGIC_VECTOR(INST_CNT_WIDTH-1 DOWNTO 0);
	SIGNAL pc_prev_q				: STD_LOGIC_VECTOR(PC_WIDTH-1 DOWNTO 0);
	SIGNAL instruction_w				: STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
	SIGNAL address_shifted2_w 		: STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
	SIGNAL zeros_helper				: STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0) := (others => '0');
BEGIN

--ROM for Instruction Memory
	inst_memory: altsyncram
	GENERIC MAP (
		operation_mode 	=> "ROM",
		width_a 			=> DATA_BUS_WIDTH,
		widthad_a 		=> ITCM_ADDR_WIDTH,
		numwords_a 	=> WORDS_NUM,
		lpm_hint 		=> "ENABLE_RUNTIME_MOD = YES,INSTANCE_NAME = ITCM",
		lpm_type 		=> "altsyncram",
		outdata_reg_a 	=> "UNREGISTERED",
		init_file 			=> "C:\intelFPGA\myWorkspace\MIPS Based MCU\Software Test Samples\Interrupt based IO\test1\bin\M9K\ITCM.hex",
		intended_device_family => "Cyclone"
	)
	PORT MAP (
		clock0 		=> clk_i,
		address_a 	=> itcm_addr_w,
		q_a 		=> instruction_w
	);
	
	-- Instructions always start on word address - not byte
	pc_q(1 DOWNTO 0) 	<= "00";
	
	-- send address to inst. memory
	G1: 
	if (WORD_GRANULARITY = True) generate -- i.e. each WORD has unique address
		itcm_addr_w <= next_pc_with_interrupts_w;
	elsif (WORD_GRANULARITY = False) generate -- i.e. each BYTE has unique address
		itcm_addr_w <= next_pc_with_interrupts_w & "00";
	end generate;
	
	-- Adder to increment PC by 4
	pc_plus4_r(1 DOWNTO 0) <= "00";
    pc_plus4_r(PC_WIDTH-1 DOWNTO 2) <= pc_q(PC_WIDTH-1 DOWNTO 2) + 1;
	
	-- Mux to select Branch Address or PC + 4        
	------------------------------------------------------------------------------------				
	next_pc_mux1_w 	<= (others => '0') WHEN rst_flag_q = '1' ELSE
					add_result_i WHEN ((Branch_ctrl_i = "10") AND (zero_i = '1')) OR ((Branch_ctrl_i = "01") AND (zero_i = '0')) ELSE -- Branch_ctrl_i = "10" -> beq, Branch_ctrl_i = "01" -> bne
					pc_plus4_r(PC_WIDTH-1 DOWNTO 2);
	-------------------------------------------------------------------------------------
	-- Mux to select Jump Address or (Branch / PC + 4)        
	------------------------------------------------------------------------------------				
	next_pc_mux2_w  <= (others => '0') WHEN rst_flag_q = '1' ELSE -- next pc address if there were no interrupts
					address_shifted2_w(PC_WIDTH-1 DOWNTO 2) WHEN Jump_ctrl_i = "11" OR Jump_ctrl_i = "10" ELSE -- jump / Jal
					alu_res_i(PC_WIDTH-1 DOWNTO 2) WHEN Jump_ctrl_i = "01" ELSE -- jr
					next_pc_mux1_w;-- no jump
					
	-- next pc if there was no interrupt - for storage in $k1
	next_pc_no_INT_o <= zeros_helper(DATA_BUS_WIDTH-1 DOWNTO PC_WIDTH) & next_pc_mux2_w & b"00";
	-- next pc if there was an interrupt
	next_pc_with_interrupts_w <= ISR_addr_i(PC_WIDTH-1 DOWNTO 2) WHEN jump_PC_to_ISR_i = '1' ELSE -- jal to ISR (so need to set PC = ISR_addr)
							next_pc_mux2_w;
	-------------------------------------------------------------------------------------
	process (clk_i)
	BEGIN
		IF(clk_i'EVENT  AND clk_i='1') THEN
			rst_flag_q <= rst_i;
		end if;
	end process;
	-------------------------------------------------------------------------------------
	PROCESS (clk_i, rst_i)
	BEGIN
		IF rst_i = '1' THEN
			pc_q(PC_WIDTH-1 DOWNTO 2) <= (OTHERS => '0') ; 
		ELSIF(clk_i'EVENT  AND clk_i='1') THEN
			pc_q(PC_WIDTH-1 DOWNTO 2) <= next_pc_with_interrupts_w;
		END IF;
	END PROCESS;
---------------------------------------------------------------------------------------
--						IPC - instruction counter register
---------------------------------------------------------------------------------------
process (clk_i , rst_i)
begin
	if rst_i = '1' then
		pc_prev_q <= (others	=> '0');
	elsif falling_edge(clk_i) then
		pc_prev_q <= pc_q;
	end if;
end process;
---------------------------------------------------------------------------------------
process (clk_i , rst_i)
begin
	if rst_i = '1' then
		inst_cnt_q <= (others => '0');
	elsif rising_edge(clk_i) then
		if pc_prev_q = pc_q then
			inst_cnt_q <= inst_cnt_q + '1';
		end if;
	end if;
end process;
---------------------------------------------------------------------------------------
	-- copy output signals - allows read inside module
	pc_o 				<= 	pc_q;
	pc_plus4_o 			<= 	pc_plus4_r;
	inst_cnt_o			<=	inst_cnt_q;
	instruction_o 		<= instruction_w;
	address_shifted2_w 	<= instruction_w(DATA_BUS_WIDTH-3 DOWNTO 0) & b"00";
END behavior;


